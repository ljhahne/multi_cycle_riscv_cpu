`ifndef IMMSRC
`define IMMSRC

`define IMMSRC_I 3'b000
`define IMMSRC_S 3'b001
`define IMMSRC_B 3'b010
`define IMMSRC_J 3'b011
`define IMMSRC_U 3'b100

`endif