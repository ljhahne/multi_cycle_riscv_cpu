`ifndef ALU
`define ALU

`define ALU_ADD 3'b000
`define ALU_SUB 3'b001
`define ALU_AND 3'b010
`define ALU_OR  3'b011
`define ALU_SLT 3'b101
`define ALU_SLL 3'b110
`define ALU_LUI 3'b100
`define ALU_DEFAULT 32'bx

`endif