`ifndef FSM
`define FSM


`define FETCH_ADRSRC 1'b0
`define FETCH_IRWRITE 1'b1
`define FETCH_ALUSRCA 2'b00
`define FETCH_ALUSRCB 2'b10
`define FETCH_ALUOP 2'b00
`define FETCH_RESULTSRC 2'b10
`define FETCH_PCUPDATE 1'b1


`define DECODE_ALUSRCA 2'b01
`define DECODE_ALUSRCB 2'b01
`define DECODE_ALUOP 2'b00


`define MEMADR_ALUSRCA 2'b10
`define MEMADR_ALUSRCB 2'b01
`define MEMADR_ALUOP 2'b00

`define EXECUTER_ALUSRCA 2'b10
`define EXECUTER_ALUSRCB 2'b00
`define EXECUTER_ALUOP 2'b10

`define EXECUTEL_ALUSRCA 2'b10
`define EXECUTEL_ALUSRCB 2'b01
`define EXECUTEL_ALUOP 2'b10


`define JAL_ALUSRCA 2'b01
`define JAL_ALUSRCB 2'b10
`define JAL_RESULTSRC 2'b00
`define JAL_ALUOP 2'b00
`define JAL_PCUPDATE 1'b1

`define BEQ_ALUSRCA 2'b10
`define BEQ_ALUSRCB 2'b00
`define BEQ_ALUOP 2'b01
`define BEQ_RESULTSRC 2'b00
`define BEQ_BRANCH 1'b1

`define MEMREAD_RESULTSRC 2'b00
`define MEMREAD_ADRSRC 1'b1

`define MEMWRITE_RESULTSRC 2'b00
`define MEMWRITE_ADRSRC 1'b1
`define MEMWRITE_MEMWRITE 1'b1

`define ALUWB_RESULTSRC 2'b00
`define ALUWB_REGWRITE 1'b1

`define MEMWB_RESULTSRC 2'b01
`define MEMWB_REGWRITE 1'b1

`define LUI_ALUSRCB 2'b01
`define LUI_ALUOP 2'b11

`define DEFAULT_ALUSRCA 2'b00
`define DEFAULT_ALUSRCB 2'b00
`define DEFAULT_RESULTSRC 2'b00
`define DEFAULT_ADRSRC 1'b0
`define DEFAULT_IRWRITE 1'b0
`define DEFAULT_ALUOP 2'b00
`define DEFAULT_PCUPDATE 1'b0
`define DEFAULT_REGWRITE 1'b0
`define DEFAULT_MEMWRITE 1'b0
`define DEFAULT_BRANCH 1'b0


`endif